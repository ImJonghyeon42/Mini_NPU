`timescale 1ns/1ps
module top_controller(
	input logic clk,
	input logic rst,
	input logic start,
	input logic [7:0] rx_data,
	input logic  rx_valid,
	output logic [7:0] tx_data, // 차선 중심 위치 (0~29)
	output logic [7:0] confidence, //신뢰도 (최대값 크기)
	output logic done_signal
);

	logic start_signal;
	logic conv_engine_done;
	logic signed [17:0] max_val_reg;
	logic [7:0] max_position_reg;
	logic [5:0]  count;
	logic [255:0] flattened_pixel_data;
	logic [7:0] pixel_row_data [0:31];
	logic signed [17:0] result_data [0:29];
	
	enum logic [2:0] {IDLE, RECEIVE_DATA, COMPUTE, FIND_MAX, SEND_RESULT} state;
	
	always_comb begin
		for( int i=0;i<32;i++) flattened_pixel_data[i*8 +: 8] = pixel_row_data[i];
	end
	
	conv_engine U0(
		.clk, .rst,
		.start(start_signal),
		.pixel_row_data(flattened_pixel_data),
		.done_signal(conv_engine_done),
		.result_data
	);

	always_ff@(posedge clk) begin
		if(rst) begin
			max_val_reg <= '0;
			state <= IDLE;
			count <= '0;
			start_signal <= '0;
			done_signal <= '0;
			tx_data <= '0;
			pixel_row_data <= '{default: '0};
			confidence <= '0;
		end
		else begin
			start_signal <= '0;
			done_signal <= 0;
			case(state) 
				IDLE : begin
				    if(start) begin 
				        state <= RECEIVE_DATA;
				        count <= '0;
				    end
				end
				RECEIVE_DATA : begin
					if(rx_valid) begin
						pixel_row_data[count[4:0]] <= rx_data;
						if(count[4:0] == 5'd31) begin
							state <= COMPUTE;
							count <= '0;
							start_signal <= '1;
						end
						else count <= count +6'd1;
					end
				end
				COMPUTE : begin
					if(conv_engine_done) begin
						state <= FIND_MAX;
						max_val_reg <= result_data[0];
						count <= 6'd1;
					end
				end
				FIND_MAX : begin
					if(result_data[count[4:0]] > max_val_reg) begin
					    max_val_reg <= result_data[count[4:0]];
					    max_position_reg <= count[4:0];
					end else if((-result_data[count[4:0]])> max_val_reg) begin
					   max_val_reg <= -result_data[count[4:0]];
					   max_position_reg <= count[4:0];
					end
					    					
					if(count[4:0] == 5'd29) begin
						state <= SEND_RESULT;
						count <= '0;
					end
					else count <= count + 6'd1;
				end
				SEND_RESULT: begin
					tx_data <= max_position_reg;
					if(max_val_reg > 255) confidence <= 8'd255;
					else confidence <= max_val_reg[7:0];
					
					done_signal <= 1'b1;
					state <= IDLE;
				end
			endcase
		end
	end
endmodule
	