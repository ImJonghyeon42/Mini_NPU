`timescale 1ns/1ps
module Fully_Connected_Layer(