`timescale 1ns/1ps
module Feature_Extractor_Fixed(
	input logic clk,
	input logic rst,
	input logic start_signal,
	input logic pixel_valid_in,
	input logic [7:0] pixel_in,
	output logic signed [21:0] final_result_out,
	output logic final_result_valid,
	output logic final_done_signal
);
	logic signed [21:0] conv_result;
	logic conv_valid;
	logic conv_done_signal;
	
	logic Activation_valid;
	logic signed [21:0] Activation_result;
	
	// ===== 22비트로 데이터 보존 (BRAM 사용) =====
	(* ram_style = "block" *) logic signed [21:0] conv_buffer [0:899];  // 16→22비트로 수정
	logic [9:0] buffer_addr;
	logic buffer_write_en;
	logic buffer_complete;
	
	// Max Pooling 입력 제어
	logic max_pool_start;
	logic conv_done_d1;
	logic [9:0] read_addr;
	logic reading_buffer;
	logic read_valid;
	logic signed [21:0] buffered_data;
	
	conv_engine_2d	U0(
		.clk, .rst, .start_signal, 
		.pixel_in, .pixel_valid(pixel_valid_in),
		.result_out(conv_result), .result_valid(conv_valid),
		.done_signal(conv_done_signal)
	);
	
	Activation_Function U1(
		.clk, .rst,
		.pixel_valid(conv_valid), .pixel_in(conv_result),
		.result_valid(Activation_valid), .result_out(Activation_result)
	);
	
	// ===== 개선된 버퍼 관리 (데이터 손실 방지) =====
	assign buffer_write_en = Activation_valid;
	
	always_ff @(posedge clk or negedge rst) begin
		if (!rst) begin
			buffer_addr <= 10'b0;
			buffer_complete <= 1'b0;
		end else if (buffer_write_en) begin
			// ✅ 수정: 22비트 전체 저장 (데이터 손실 없음)
			conv_buffer[buffer_addr] <= Activation_result;  // 전체 22비트 보존
			
			if (buffer_addr == 899) begin  // 30x30 = 900
				buffer_addr <= 10'b0;
				buffer_complete <= 1'b1;
				$display("Feature Buffer 완료: 900개 픽셀 저장됨");
			end else begin
				buffer_addr <= buffer_addr + 1;
			end
		end else if (!conv_done_signal) begin
			buffer_complete <= 1'b0;
		end
	end
	
	// Conv 완료 감지
	always_ff @(posedge clk or negedge rst) begin
		if (!rst) begin
			conv_done_d1 <= 1'b0;
		end else begin
			conv_done_d1 <= conv_done_signal;
		end
	end
	
	assign max_pool_start = buffer_complete && !conv_done_d1;
	
	// ===== 개선된 버퍼 읽기 =====
	always_ff @(posedge clk or negedge rst) begin
		if (!rst) begin
			read_addr <= 10'b0;
			reading_buffer <= 1'b0;
			read_valid <= 1'b0;
		end else if (max_pool_start) begin
			reading_buffer <= 1'b1;
			read_addr <= 10'b0;
			read_valid <= 1'b1;
			$display("Max Pooling 시작: 900개 픽셀 처리");
		end else if (reading_buffer) begin
			if (read_addr == 899) begin
				read_addr <= 10'b0;
				reading_buffer <= 1'b0;
				read_valid <= 1'b0;
				$display("버퍼 읽기 완료");
			end else begin
				read_addr <= read_addr + 1;
			end
		end
	end
	
	// ✅ 수정: 22비트 데이터 그대로 사용 (부호 확장 불필요)
	assign buffered_data = conv_buffer[read_addr];
	
	Max_Pooling #( .IMG_WIDTH(30), .IMG_HEIGHT(30))
	U2 (
		.clk, .rst, 
		.start_signal(max_pool_start),
		.pixel_in(buffered_data), 
		.pixel_valid(read_valid),
		.result_out(final_result_out), 
		.result_valid(final_result_valid), 
		.done_signal(final_done_signal)
	);
	
endmodule